module CDAC_13_11 (
	inout[5:0]  CB,
	inout CT,
	inout  VSS,
 	inout VDD,
	inout  VNW,
 	inout VPW
);

wire AVDD;
wire AVSS;
wire [9:0] CBC;
MOM2D I_0_1 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_0_2 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_0_3 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_0_4 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_0_5 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_0_6 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_0_7 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_0_8 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_0_9 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_0_10 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
SC7P5T_INVX1_SSC14R  I_1_0(.Z(CBC[9]), .A(CB[5]), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_1_1 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_1_2 ( .CB(CBC[9]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_1_3 ( .CB(CBC[9]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_1_4 ( .CB(CBC[9]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_1_5 ( .CB(CBC[9]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_1_6 ( .CB(CBC[9]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_1_7 ( .CB(CBC[9]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_1_8 ( .CB(CBC[9]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_1_9 ( .CB(CBC[9]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_1_10 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
SC7P5T_INVX1_SSC14R  I_2_0(.Z(CBC[8]), .A(CB[4]), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_2_1 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_2_2 ( .CB(CBC[8]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_2_3 ( .CB(CBC[8]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_2_4 ( .CB(CBC[8]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_2_5 ( .CB(CBC[8]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_2_6 ( .CB(CBC[8]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_2_7 ( .CB(CBC[8]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_2_8 ( .CB(CBC[8]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_2_9 ( .CB(CBC[8]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_2_10 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
SC7P5T_INVX1_SSC14R  I_3_0(.Z(CBC[7]), .A(CB[5]), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_3_1 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_3_2 ( .CB(CBC[7]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_3_3 ( .CB(CBC[7]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_3_4 ( .CB(CBC[7]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_3_5 ( .CB(CBC[7]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_3_6 ( .CB(CBC[7]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_3_7 ( .CB(CBC[7]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_3_8 ( .CB(CBC[7]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_3_9 ( .CB(CBC[7]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_3_10 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
SC7P5T_INVX1_SSC14R  I_4_0(.Z(CBC[6]), .A(CB[3]), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_4_1 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_4_2 ( .CB(CBC[6]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_4_3 ( .CB(CBC[6]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_4_4 ( .CB(CBC[6]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_4_5 ( .CB(CBC[6]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_4_6 ( .CB(CBC[6]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_4_7 ( .CB(CBC[6]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_4_8 ( .CB(CBC[6]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_4_9 ( .CB(CBC[6]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_4_10 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
SC7P5T_INVX1_SSC14R  I_5_0(.Z(CBC[5]), .A(CB[5]), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_5_1 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_5_2 ( .CB(CBC[5]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_5_3 ( .CB(CBC[5]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_5_4 ( .CB(CBC[5]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_5_5 ( .CB(CBC[5]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_5_6 ( .CB(CBC[5]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_5_7 ( .CB(CBC[5]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_5_8 ( .CB(CBC[5]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_5_9 ( .CB(CBC[5]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_5_10 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
SC7P5T_INVX1_SSC14R  I_6_0(.Z(CBC[4]), .A(CB[4]), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_6_1 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_6_2 ( .CB(CBC[4]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_6_3 ( .CB(CBC[4]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_6_4 ( .CB(CBC[4]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_6_5 ( .CB(CBC[4]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_6_6 ( .CB(CBC[4]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_6_7 ( .CB(CBC[4]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_6_8 ( .CB(CBC[4]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_6_9 ( .CB(CBC[4]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_6_10 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
SC7P5T_INVX1_SSC14R  I_7_0(.Z(CBC[3]), .A(CB[5]), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_7_1 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_7_2 ( .CB(CBC[3]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_7_3 ( .CB(CBC[3]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_7_4 ( .CB(CBC[3]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_7_5 ( .CB(CBC[3]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_7_6 ( .CB(CBC[3]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_7_7 ( .CB(CBC[3]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_7_8 ( .CB(CBC[3]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_7_9 ( .CB(CBC[3]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_7_10 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
SC7P5T_INVX1_SSC14R  I_8_0(.Z(CBC[2]), .A(CB[2]), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_8_1 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_8_2 ( .CB(CBC[2]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_8_3 ( .CB(CBC[2]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_8_4 ( .CB(CBC[2]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_8_5 ( .CB(CBC[2]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_8_6 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_8_7 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_8_8 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_8_9 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_8_10 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
SC7P5T_INVX1_SSC14R  I_9_0(.Z(CBC[1]), .A(CB[1]), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_9_1 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_9_2 ( .CB(CBC[1]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_9_3 ( .CB(CBC[1]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_9_4 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_9_5 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_9_6 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_9_7 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_9_8 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_9_9 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_9_10 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
SC7P5T_INVX1_SSC14R  I_10_0(.Z(CBC[0]), .A(CB[0]), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_10_1 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_10_2 ( .CB(CBC[0]), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_10_3 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_10_4 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_10_5 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_10_6 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_10_7 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_10_8 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_10_9 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_10_10 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_11_1 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2 I_11_2 ( .CB(VSS), .CT(CT), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_11_3 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_11_4 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_11_5 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_11_6 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_11_7 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_11_8 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_11_9 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_11_10 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_12_1 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_12_2 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_12_3 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_12_4 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_12_5 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_12_6 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_12_7 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_12_8 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_12_9 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
MOM2D I_12_10 ( .CB(VSS), .CT(VSS), .VDD(VDD), .VSS(VSS), .VPW(VPW), .VNW(VNW));
endmodule

